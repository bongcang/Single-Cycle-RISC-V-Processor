`timescale 1ns / 1ps

module processor (
    input clk, reset,
    
    output [31:0] Result
    );
    
endmodule
